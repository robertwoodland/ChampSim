import *TO_SUBSTITUTE_FILE*::*;
import BrPred::*;

export mkDirPredictor;
export DirPredTrainInfo(..);

module mkDirPredictor(DirPredictor#(DirPredTrainInfo));
    let m <- *TO_SUBSTITUTE_MODULE*;
    return m;
endmodule