typedef 128 GlobalHistoryLength;
typedef 8 MaxSpecSize;
