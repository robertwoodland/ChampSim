typedef 128 GlobalHistoryLength;