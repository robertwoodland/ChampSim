typedef 64 AddrSz;
typedef Bit#(AddrSz) Addr;
typedef 1 SupSize;
typedef Bit#(TLog#(TAdd#(SupSize, 1))) SupCnt;